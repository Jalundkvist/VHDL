package car_state_pkg is

type car_state_t is (parked, is_driving, ignition_on);

end package;