library IEEE;
use IEEE.std_logic_1164.all;

ENTITY 7seg is
	port
	(
	input : in std_logic_vector; (3 downto 0);
	output : out std_logic_vector ( 6 downto 0)
	);
end 7seg;

architecture 7seg of 7seg is
	begin
	
	
end architecture;